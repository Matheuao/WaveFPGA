library ieee;
use ieee.numeric_std.all;

package vector_types is
  type signed_vector is array (natural range <>) of signed;
  
end package vector_types;


package body vector_types is
end package body vector_types;
