library ieee;
use ieee.std_logic_1164.all;

package dwt_types is

  -- Versões da transformada DWT
  type dwt_transform_version is (
    DWT_V1,
    DWT_V2
    -- NDWT_V3, etc.
  );

end package dwt_types;

package body dwt_types is
end package body dwt_types;
