library ieee;
use ieee.std_logic_1164.all;

package ndwt_types is

  -- Versões da transformada NDWT
  type ndwt_transform_version is (
    NDWT_V1,
    NDWT_V2
    -- NDWT_V3, etc.
  );

end package ndwt_types;

package body ndwt_types is
end package body ndwt_types;
